while (free_time) begin
	$display ("Work on 385");
end