always begin
	#5 clk = ~clk;
end

//#5 delays execution by 5 time units