for (i=0; i < 16; i = i + 1) begin
	$display("Current value of i is %d", i);
end