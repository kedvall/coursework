case(address)
	0 : $display ("It is 12:00");
	1 : $display ("Need sleep...");
	2 : $display ("Help meeee");
	default : $display ("Must finish this");
endcase