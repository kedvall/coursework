repeat (16) begin //Repeats code block 16 times
	$display("Current value of i is %d", i);
	i = i+1;
end