initial begin //For use in testbench ONLY
	clk = 0;
	reset = 0'
	req = 0;
end 